library ieee;
use ieee.std_logic_1164.all;

entity seven_segments is

	port(
	sw : in std_logic_vector(2 downto 0);
	pb: in std_logic;
	hex0: out std_logic_vector(0 to 7));
end seven_segments;

architecture seven_segment_arch of seven_segments is
	begin
		with pb & sw select
		hex0 <= "00000011" when "0000", --0
				"10011111" when "0001", --1
				"00100101" when "0010", --2
				"00001101" when "0011", --3
				"10011001" when "0100", --4
				"01001001" when "0101", --5
				"01000001" when "0110", --6
				"00011111" when "0111", --7
				"00000001" when "1000", --8
				"00011001" when "1001", --9
				"00010001" when "1010", --A
				"11000001" when "1011", --b
				"01100011" when "1100", --C
				"10000101" when "1101", --d
				"01100001" when "1110", --E
				"01110001" when "1111", --F
				"11111111" when others;
end seven_segment_arch;